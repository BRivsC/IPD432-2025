// Módulo top pregunta 3 tarea 1
// Incluye un debouncer y una máquina de estados PB_FSM de tipo Moore
module T1_design1 #(
    parameter N_DEBOUNCER_DELAY = 10,
    parameter N_INCREMENT_DELAY_CONTINUOUS = 5
)(
    input   logic   clk,
    input   logic   resetN,
    input   logic   PushButton,
    output  logic   IncPulse_out
);

endmodule